library verilog;
use verilog.vl_types.all;
entity lab02_vlg_check_tst is
    port(
        output_1        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab02_vlg_check_tst;
