library verilog;
use verilog.vl_types.all;
entity part2 is
    port(
        D               : out    vl_logic;
        A               : in     vl_logic;
        B               : in     vl_logic;
        C               : in     vl_logic
    );
end part2;
