library verilog;
use verilog.vl_types.all;
entity lab04_vlg_check_tst is
    port(
        OUT_GNT0        : in     vl_logic;
        OUT_GNT1        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end lab04_vlg_check_tst;
